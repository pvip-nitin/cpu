		mem[16'hFFFF] <= 16'h10;
		mem[16'hFFFE] <= 16'h20;
		mem[16'hFFFD] <= 16'h30;
