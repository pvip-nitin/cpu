module cpu_top
  #(
    ADDR_WIDTH = 16,
    DATA_WIDTH = 16
    )
   (
     cr_if      crIf,
     read_if    instrIf,
     read_if    rdataIf,
     write_if   wdataIf
    );


endmodule
