interface cr_if
(
  input     clk,
  input     rstn
);

endinterface
